parameter OFF = 8'b11111111;
parameter N0  = 8'b11000000;
parameter N1  = 8'b11111001;
parameter N2  = 8'b10100100;
parameter N3  = 8'b10110000;
parameter N4  = 8'b10011001;
parameter N5  = 8'b10010010;
parameter N6  = 8'b10000010;
parameter N7  = 8'b11111000;
parameter N8  = 8'b10000000;
parameter N9  = 8'b10011000;
parameter A   = 8'b10001000;
parameter C   = 8'b11000110;
parameter E   = 8'b10000110;
parameter G   = 8'b11000010;
parameter H   = 8'b10001001;
parameter I   = 8'b11001111;
parameter J   = 8'b11100001;
parameter K   = 8'b10001010;
parameter L   = 8'b11000111;
parameter M   = 8'b11101010;
parameter N   = 8'b10101011;
parameter O   = 8'b10100011;
parameter P   = 8'b10001100;
parameter R   = 8'b11001100;
parameter S   = 8'b10010010;
parameter T   = 8'b10000111;
parameter U   = 8'b11000001;
parameter Y   = 8'b10010001;
